* Author: L. Schindler
* Version: 1.5.1
* Last modification date: 18 June 2020
* Last modification by: L. Schindler

* Copyright (c) 2018-2020 Lieze Schindler, Stellenbosch University

* Permission is hereby granted, free of charge, to any person obtaining a copy
* of this cell library and associated documentation files (the "Library"), to deal
* in the Library without restriction, including without limitation the rights
* to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
* copies of the Library, and to permit persons to whom the Library is
* furnished to do so, subject to the following conditions:

* The above copyright notice and this permission notice shall be included in all
* copies or substantial portions of the Library.

* THE LIBRARY IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
* IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
* FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
* AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
* LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
* OUT OF OR IN CONNECTION WITH THE LIBRARY OR THE USE OR OTHER DEALINGS IN THE
* LIBRARY.

*For questions about the library, contact Lieze Schindler, 17528283@sun.ac.za

*$Ports 			  a q
.subckt LSMITLL_JTLT a q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.2p
.param ICreceive=1.6
.param ICtrans=2.5
.param Lptl=2p
.param LB=2p
.param BiasCoef=0.7
.param RD=1.36
.param B1=ICreceive
.param B2=ICtrans/1.25
.param B3=ICtrans
.param IB1=B1*Ic0*BiasCoef
.param IB2=(B2+B3)*Ic0*BiasCoef
.param L1=Lptl
.param L2=Phi0/(2*B1*Ic0)
.param L3=(Phi0/(2*B2*Ic0))/2
.param L4=L3
.param L5=Lptl
.param LP1=LP
.param LP2=LP
.param LP3=LP
.param LB1=LB
.param LB2=LB
.param RB1=B0Rs/B1   
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet+LP
.param LRB3=(RB3/Rsheet)*Lsheet+LP
B1         6          7          jjmit area=B1
B2         9          10         jjmit area=B2
B3         12         13         jjmit area=B3
IB1         0          18        pwl(0      0 5p IB1)
IB2         0          19        pwl(0      0 5p IB2)
L1         a          6          L1        
L2         6          9          L2     
L3         9          16         L3       
L4         16         12         L4        
L5         12         17         L5        
LB1        6          18         LB1        
LB2        16         19         LB2        
LP1        0          7          LP1      
LP2        0          10         LP2      
LP3        0          13         LP3
LRB1       0          8          LRB1     
LRB2       0          11         LRB2     
LRB3       0          14         LRB3    
RB1        8          6          RB1     
RB2        11         9          RB2    
RB3        14         12         RB3     
RD         17         q          RD              
.ends